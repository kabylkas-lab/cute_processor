// -----------------------------------------------------------------------------
// Register
// -----------------------------------------------------------------------------
module regn(
    // -------------------------------------------------------------------------
    // Inputs
    // -------------------------------------------------------------------------
    input wire clk,
    input wire enable,
    input wire signed [8:0] a0,
    // -------------------------------------------------------------------------
    
    // Register
    output reg signed [8:0] reg0
    // -------------------------------------------------------------------------
);

// -----------------------------------------------------------------------------
// Register update
// -----------------------------------------------------------------------------
always@ (posedge clk) begin
    if (enable) reg0 <= a0;
end
// -----------------------------------------------------------------------------
endmodule