// -----------------------------------------------------------------------------
// Register
// -----------------------------------------------------------------------------
module regn(
    // -------------------------------------------------------------------------
    // Inputs
    // -------------------------------------------------------------------------
    input wire clk,
    input wire Reset,
    input wire [8:0] a0,
    // -------------------------------------------------------------------------
    
    // Register
    output reg reg0
    // -------------------------------------------------------------------------
);

// -----------------------------------------------------------------------------
// Register update
// -----------------------------------------------------------------------------
always@ (posedge clk) begin
    if (Reset) reg0 = 9d0;
    else reg0 = a0;
end
// -----------------------------------------------------------------------------

endcase
// -----------------------------------------------------------------------------
